LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEM_A_READ_COUNTER IS  
	PORT(CLK, RST, EN: IN STD_LOGIC;
	ADDR_B: IN UNSIGNED(9 DOWNTO 0);                    -- EN IS RD_A FROM CONTROL UNIT, ADDR_B IS THE ADDRESS OF B MEMORY USED AS MASK
	ADDR: OUT UNSIGNED(9 DOWNTO 0));
END MEM_A_READ_COUNTER;

ARCHITECTURE behavior OF MEM_A_READ_COUNTER IS
SIGNAL ADDR_AUX : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";


BEGIN
PROCESS(CLK, RST)
BEGIN
	IF RST = '1' THEN
		ADDR_AUX <= (OTHERS => '0');  -- ASYNC RESET
	ELSE 
		IF (CLK = '1' AND CLK'EVENT) THEN
			IF EN = '1' THEN
				ADDR_AUX <= STD_LOGIC_VECTOR(UNSIGNED(ADDR_AUX) + 1);	
			ELSE
				ADDR_AUX <= STD_LOGIC_VECTOR(UNSIGNED(ADDR_AUX));
			END IF;
		END IF;
	END IF;
END PROCESS;

ADDR <= ADDR_B - UNSIGNED(ADDR_AUX);

END behavior;
		
	