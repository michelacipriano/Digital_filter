LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEMORY_A IS
	PORT (ADDRESS_M_A: IN UNSIGNED(9 DOWNTO 0);
	      UNDERFLOW: IN STD_LOGIC;
	      DATA_IN_M: IN SIGNED(7 DOWNTO 0); 
	      CS_M_A,WR_M_A,RD_M_A,CLK_A: IN STD_LOGIC;
	       Q_OUT: OUT SIGNED (7 DOWNTO 0));
END MEMORY_A;

ARCHITECTURE BEHAVIOR OF MEMORY_A IS

TYPE MAT IS ARRAY (1023 DOWNTO 0) OF SIGNED(7 DOWNTO 0); --1023 CAMPIONI, CIASCUNO DEI QUALI E' UN VETTORE DA 8 BIT
SIGNAL MEMORY_SIG: MAT;
BEGIN
P0: PROCESS(CLK_A)  --PROCESS CHE, PER OGNI CICLO DI CLK, INSERISCE OGNI VETTORE DI 8 BIT "DATA_IN" IN INGRESSO NELL'ELEMENTO DI MATRICE DI POSTO "ADDRESS"
BEGIN
	IF (CLK_A = '1' AND CLK_A'EVENT) THEN
		IF CS_M_A = '1' AND WR_M_A = '1' THEN
			MEMORY_SIG(TO_INTEGER(ADDRESS_M_A)) <= DATA_IN_M;
		END IF;
	END IF;

END PROCESS P0;

P1: PROCESS(ADDRESS_M_A) --PROCESS CHE, IN MANIERA ASINCRONA, LEGGE IL VETTORE DI 8 BIT NELL'ELEMENTO DI MATRICE DI POSTO "ADDRESS" E LO MANDA IN OUTPUT
	BEGIN
		IF CS_M_A = '1' AND RD_M_A = '1' AND UNDERFLOW = '0' THEN
			Q_OUT <= MEMORY_SIG(TO_INTEGER(ADDRESS_M_A));
		ELSE
			Q_OUT <= (OTHERS => '0');
		END IF;

END PROCESS P1;


END BEHAVIOR;