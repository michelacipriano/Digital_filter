LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY MEMORY_B IS
	PORT (ADDRESS_M_B: IN UNSIGNED(9 DOWNTO 0);
	      DATA_OUT: IN SIGNED(7 DOWNTO 0); 
	      CS_M_B,WR_M_B,CLK_B: IN STD_LOGIC);
END MEMORY_B;

ARCHITECTURE BEH OF MEMORY_B IS
TYPE MAT IS ARRAY (1023 DOWNTO 0) OF SIGNED(7 DOWNTO 0);
SIGNAL MEMORY_SIG: MAT;
BEGIN

P0: PROCESS(CLK_B)  
BEGIN
	IF (CLK_B = '1' AND CLK_B'EVENT) THEN
		IF CS_M_B = '1' AND WR_M_B = '1' THEN
			MEMORY_SIG(TO_INTEGER(ADDRESS_M_B)) <= DATA_OUT;
		ELSE
			MEMORY_SIG(TO_INTEGER(ADDRESS_M_B)) <= MEMORY_SIG(TO_INTEGER(ADDRESS_M_B));
		END IF;
	END IF;

END PROCESS P0;
END BEH;
