LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY filtering_function IS
PORT(X : IN SIGNED (7 DOWNTO 0);
     INV: IN SIGNED(0 DOWNTO 0);
     LD, SH: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
     LOC: IN NATURAL;
     CLOCK, RESET, D, RST_SUM : IN STD_LOGIC;
     Y : OUT SIGNED (10 DOWNTO 0));
END filtering_function;


ARCHITECTURE behavior OF filtering_function IS

SIGNAL ADD_LOAD1, ADD_MUX, ADD_XOR, ADD_SHIFTED, X_EXT, INV_EXT, PARTIAL_SUM, SUM_BUFFER_MUX, SUM_BUFFER : SIGNED (10 DOWNTO 0) := (OTHERS => '0');
SIGNAL SEL: STD_LOGIC := '0';

COMPONENT ADDER IS 
	PORT (a, b : IN SIGNED(10 DOWNTO 0);
     	 carry_in: SIGNED;
      	 final_sum: OUT SIGNED(10 downto 0));
END COMPONENT;

COMPONENT generic_reg is
	PORT( D: IN SIGNED(10 DOWNTO 0);
	      LD, SH, CLOCK, RESET: IN STD_LOGIC;
	      N : IN NATURAL;
	      Q: OUT SIGNED(10 DOWNTO 0));
END COMPONENT;

COMPONENT  D_flip_flop is
	PORT ( D, CLK, CL: IN STD_LOGIC;
		Q: OUT STD_LOGIC);
end COMPONENT;

COMPONENT mux2 IS
	PORT(a, b : IN SIGNED(10 DOWNTO 0);
	inv : IN STD_LOGIC;
	c : OUT SIGNED (10 DOWNTO 0));
END COMPONENT;

COMPONENT EXTENDER IS 
	PORT(data : IN SIGNED (7 DOWNTO 0);
	extended_data : OUT SIGNED (10 DOWNTO 0));
END COMPONENT;


BEGIN
INV_EXT <= resize(inv,inv_ext'length);

EXT: EXTENDER PORT MAP(X, X_EXT); 

SHIFTER : GENERIC_REG PORT MAP(X_EXT, LD(0), SH(0), CLOCK, RESET, LOC, ADD_SHIFTED); 

LOAD1 : GENERIC_REG PORT MAP(ADD_SHIFTED, LD(1), SH(1), CLOCK, RESET, LOC, ADD_LOAD1);

ADD_XOR <= ADD_LOAD1 XOR INV_EXT;

ADD : ADDER  PORT MAP (ADD_MUX, SUM_BUFFER_MUX, INV, PARTIAL_SUM);

LOAD2 : GENERIC_REG PORT MAP(PARTIAL_SUM, LD(2), SH(2), CLOCK, RESET, LOC, SUM_BUFFER);

DFF: D_FLIP_FLOP PORT MAP(D,CLOCK, RESET, SEL);

MUX_SUM1: MUX2 PORT MAP( ADD_XOR, "00000000000", SEL, ADD_MUX);
MUX_SUM_F: MUX2 PORT MAP( SUM_BUFFER, "00000000000", RST_SUM, SUM_BUFFER_MUX);


Y <= SUM_BUFFER;


END behavior;

     
