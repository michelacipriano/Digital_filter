LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEM_B_WR_COUNTER IS
	PORT(CLK, RST, EN, DONE: IN STD_LOGIC;  --EN IS WR_B, ACTIVATED IN WRITING_B_STATUS IN THE CU
        ADDR: OUT UNSIGNED(9 DOWNTO 0));	-- DONE IS THE TERMINAL COUNT, ACTIVATED IN DONE_STATE IN THE CU
END MEM_B_WR_COUNTER;

ARCHITECTURE behavior OF MEM_B_WR_COUNTER IS

SIGNAL ADDR_OUT : STD_LOGIC_VECTOR(9 DOWNTO 0):= (OTHERS => '0');
BEGIN
PROCESS(CLK, RST)
BEGIN
	IF RST = '1' THEN               -- ASYNCHRONOUS RESET
		ADDR_OUT <= (OTHERS => '0');
	ELSE 
		IF (CLK = '1' AND CLK'EVENT) THEN
			IF (EN = '1' AND DONE = '0') THEN
				   ADDR_OUT <= STD_LOGIC_VECTOR(UNSIGNED(ADDR_OUT) + 1);	
			ELSE
				   ADDR_OUT <= STD_LOGIC_VECTOR(UNSIGNED(ADDR_OUT));	
			END IF;
		END IF;		
	END IF;

END PROCESS;
ADDR <= UNSIGNED(ADDR_OUT);
END behavior;
		
	