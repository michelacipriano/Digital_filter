LIBRARY IEEE;
USE ieee.std_logic_1164.all;       -- CHECKED AND APPROVED ;-)
USE IEEE.NUMERIC_STD.ALL;

ENTITY MEM_A_WR_COUNTER IS
	PORT(CLK, RST, EN, START: IN STD_LOGIC;                           -- EN IS WR_A, CONTROLLED BY CU;  RESET ASYNCHRONOUS
	ADDR: OUT UNSIGNED(9 DOWNTO 0);			           -- MEMORY_HAS_WRITTEN <= '1' --> LET THE CU PASS TO THE NEXT STATE
	MEM_A_HAS_WRITTEN_M : OUT STD_LOGIC);
END MEM_A_WR_COUNTER;

ARCHITECTURE behavior OF MEM_A_WR_COUNTER IS
SIGNAL ADDR_AUX: STD_LOGIC_VECTOR(9 DOWNTO 0) := "0000000000";
SIGNAL MEMORY_HAS_WRITTEN_AUX: STD_LOGIC;

BEGIN
PROCESS(CLK, RST)
BEGIN
	
	IF RST = '1' THEN
		ADDR_AUX <= "0000000000";
		MEMORY_HAS_WRITTEN_AUX <= '0';
	ELSIF (CLK = '1' AND CLK'EVENT) THEN
	 	IF EN = '1' THEN
			IF (ADDR_AUX = "1111111111") THEN
 			        ADDR_AUX <= ADDR_AUX;
				MEMORY_HAS_WRITTEN_AUX <= '1';
			ELSE
				ADDR_AUX <= STD_LOGIC_VECTOR(UNSIGNED(ADDR_AUX) + 1);
				MEMORY_HAS_WRITTEN_AUX <= '0';
			END IF;
		 ELSE
			ADDR_AUX <= ADDR_AUX;
			MEMORY_HAS_WRITTEN_AUX <= MEMORY_HAS_WRITTEN_AUX;
		END IF;
	ELSE
		ADDR_AUX <= ADDR_AUX;
		MEMORY_HAS_WRITTEN_AUX <= MEMORY_HAS_WRITTEN_AUX;
	END IF;

END PROCESS;
ADDR <= UNSIGNED(ADDR_AUX);
MEM_A_HAS_WRITTEN_M <= MEMORY_HAS_WRITTEN_AUX;
END behavior;
		
	