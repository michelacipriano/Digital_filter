LIBRARY IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE STD.textio.all;
USE ieee.std_logic_textio.all;

ENTITY TB_GM IS
END TB_GM;

ARCHITECTURE TESTBENCH OF TB_GM IS

COMPONENT ACTIVE_FILTER_TB IS
	PORT(DATA: IN SIGNED(7 DOWNTO 0);
	     CLOCK,START: IN STD_LOGIC;
	     Y_OUT: OUT SIGNED(7 DOWNTO 0);
	     DONE: OUT STD_LOGIC);
END COMPONENT;

SIGNAL CLK_AUX : STD_LOGIC;

SIGNAL DATA_IN : SIGNED (7 DOWNTO 0) := "00000000";
SIGNAL CONTATORE : INTEGER := 0;
SIGNAL RIGHE : INTEGER := 1;

SIGNAL START_AUX : STD_LOGIC := '1';
SIGNAL DONE_AUX : STD_LOGIC := '0';
SIGNAL Y_OUT_AUX : SIGNED (7 DOWNTO 0);

SIGNAL RESTART : STD_LOGIC := '0';

BEGIN

BENCH : ACTIVE_FILTER_TB PORT MAP(DATA_IN, CLK_AUX, START_AUX, Y_OUT_AUX, DONE_AUX);

IO_BENCH : PROCESS(CLK_AUX)
VARIABLE RIGA_IN : line;
FILE dati : text IS IN "dati.txt";
VARIABLE BYTE : STD_LOGIC_VECTOR(7 DOWNTO 0);

VARIABLE RIGA_OUT : line;
FILE DATI_OUT  : text OPEN write_mode IS "dati_out.txt";
VARIABLE BYTE_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);

VARIABLE RIGA_IN2 : line;
FILE dati2 : text IS IN "dati2.txt";
VARIABLE BYTE2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
IF (CLK_AUX = '1' AND CLK_AUX'EVENT) THEN
	
        IF NOT(endfile(dati)) THEN
          	readline(dati, RIGA_IN);
          	read(RIGA_IN, BYTE);
		DATA_IN <= SIGNED(BYTE);
	END IF;

	IF CONTATORE < 1035 THEN
		CONTATORE <= CONTATORE + 1;
	ELSIF RIGHE <= 1024 THEN 
		BYTE_OUT := STD_LOGIC_VECTOR(Y_OUT_AUX);
		WRITE(RIGA_OUT, BYTE_OUT);
		WRITELINE(dati_out, RIGA_OUT);
		RIGHE <= RIGHE +1;
		CONTATORE <= 1025;
	END IF;

	IF (RESTART = '1' AND RIGHE = 1025) THEN
		IF NOT(endfile(dati2)) THEN
          		readline(dati2, RIGA_IN2);
          		read(RIGA_IN2, BYTE2);
			DATA_IN <= SIGNED(BYTE2);
		END IF;
	END IF;

END IF;
END PROCESS IO_BENCH;

CLOCKING : PROCESS
BEGIN
CLK_AUX <= '1';
WAIT FOR 50 ns;
CLK_AUX <= '0';
WAIT FOR 50 ns;
END PROCESS CLOCKING;


PREPARE_RESTART : PROCESS
BEGIN
WAIT FOR 1500 us;
START_AUX <= '0';
WAIT FOR 100 ns;
RESTART <= '1';
START_AUX <= '1';
END PROCESS PREPARE_RESTART;

END TESTBENCH;

