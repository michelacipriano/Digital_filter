LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY ACTIVE_FILTER_TB IS
	PORT(DATA: IN SIGNED(7 DOWNTO 0);
	     CLOCK,START: IN STD_LOGIC;
	     Y_OUT: OUT SIGNED(7 DOWNTO 0); --Y_OUT IS AN OUTPUT, ONLY DIFFERENCE WITH RESPECT TO THE MAIN FILE
	     DONE: OUT STD_LOGIC);
END ACTIVE_FILTER_TB;

ARCHITECTURE BEH OF ACTIVE_FILTER_TB IS
SIGNAL RESET_SIG: STD_LOGIC;
SIGNAL X_SIG, Y_SAT_SIG: SIGNED(7 DOWNTO 0);
SIGNAL WR_A_SIG, WR_B_SIG, CS_A_SIG, CS_B_SIG, RD_A_SIG, RD_B_SIG: STD_LOGIC;
SIGNAL N_SHIFT_SIG: NATURAL;
SIGNAL INV_SIG: SIGNED(0 DOWNTO 0);
SIGNAL SH_SIG, LD_SIG : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL UPDATE_ADD_SIG, DONE_SIG, D_SIG, RESET_SUM_SIG, EN_SAT_SIG: STD_LOGIC;
SIGNAL MEM_A_HAS_WRITTEN_SIG, UNDERFLOW_SIG: STD_LOGIC;
SIGNAL MEM_A_ADDRESS_SIG, MEM_B_ADDRESS_SIG: UNSIGNED(9 DOWNTO 0);

COMPONENT CU IS
	PORT( START ,MEM_A_HAS_WRITTEN, CLOCK, RESET: IN STD_LOGIC;
	WR_A, RD_A, WR_B, RD_B, CS_A, CS_B, DONE, D, UPDATE_AD, RESET_SUM, EN_SAT: OUT STD_LOGIC;
	SH, LD: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	INV: OUT SIGNED;
	N_SHIFT: OUT NATURAL);
END COMPONENT;


COMPONENT MEMORY_A IS
	PORT (ADDRESS_M_A: IN UNSIGNED(9 DOWNTO 0);
	      UNDERFLOW: IN STD_LOGIC;
	      DATA_IN_M: IN SIGNED(7 DOWNTO 0); 
	      CS_M_A,WR_M_A,RD_M_A,CLK_A: IN STD_LOGIC;
	      Q_OUT: OUT SIGNED (7 DOWNTO 0));
END COMPONENT;

COMPONENT MEMORY_B IS
	PORT (ADDRESS_M_B: IN UNSIGNED(9 DOWNTO 0);
	      DATA_OUT: IN SIGNED(7 DOWNTO 0); 
	      CS_M_B,WR_M_B,CLK_B: IN STD_LOGIC);
END COMPONENT;

COMPONENT DP IS
	PORT(X: IN SIGNED(7 DOWNTO 0);
	     CLOCK, START, RESET: IN STD_LOGIC;
	     WR_A, WR_B, CS_A, CS_B, RD_A, RD_B: IN STD_LOGIC;
	     N_SHIFT: IN NATURAL;
	     INV: IN SIGNED (0 DOWNTO 0);
	     SH, LD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	     UPDATE_ADD, DONE, D, RESET_SUM, EN_SAT: IN STD_LOGIC;
	     MEM_A_HAS_WRITTEN_DP, UNDERFLOW: OUT STD_LOGIC;
	     MEM_A_ADDRESS, MEM_B_ADDRESS: OUT UNSIGNED(9 DOWNTO 0);
	     Y_SAT: OUT SIGNED(7 DOWNTO 0));
END COMPONENT;

BEGIN

CONTROL_UNIT: CU PORT MAP(START, MEM_A_HAS_WRITTEN_SIG, CLOCK, RESET_SIG, WR_A_SIG, RD_A_SIG, WR_B_SIG, RD_B_SIG, CS_A_SIG, CS_B_SIG, 
			DONE_SIG, D_SIG, UPDATE_ADD_SIG, RESET_SUM_SIG, EN_SAT_SIG, SH_SIG, LD_SIG, INV_SIG, N_SHIFT_SIG);

MEM_A: MEMORY_A PORT MAP(MEM_A_ADDRESS_SIG, UNDERFLOW_SIG, DATA, CS_A_SIG, WR_A_SIG, RD_A_SIG, CLOCK, X_SIG);

MEM_B: MEMORY_B PORT MAP(MEM_B_ADDRESS_SIG, Y_SAT_SIG, CS_B_SIG, WR_B_SIG, CLOCK);

DATAPATH: DP PORT MAP(X_SIG, CLOCK, START, RESET_SIG, WR_A_SIG, WR_B_SIG, CS_A_SIG, CS_B_SIG, RD_A_SIG, RD_B_SIG,
			N_SHIFT_SIG, INV_SIG, SH_SIG, LD_SIG, UPDATE_ADD_SIG, DONE_SIG, D_SIG, RESET_SUM_SIG, EN_SAT_SIG,
			MEM_A_HAS_WRITTEN_SIG, UNDERFLOW_SIG, MEM_A_ADDRESS_SIG, MEM_B_ADDRESS_SIG, Y_SAT_SIG);

RESET_SIG <= '1' WHEN (START = '1' AND DONE_SIG = '1' AND START'EVENT) ELSE '0';

Y_OUT <= Y_SAT_SIG;

DONE <= DONE_SIG;

END BEH;

