LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY DP IS
	PORT(--INPUT
	     X: IN SIGNED(7 DOWNTO 0);
	     CLOCK, START, RESET: IN STD_LOGIC;
	     --CONTROL SIGNALS
	     WR_A, WR_B, CS_A, CS_B, RD_A, RD_B: IN STD_LOGIC;
	     N_SHIFT: IN NATURAL;
	     INV: IN SIGNED (0 DOWNTO 0);
	     SH, LD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	     UPDATE_ADD, DONE, D, RESET_SUM, EN_SAT: IN STD_LOGIC;
	     --STATUS SIGNALS
	     MEM_A_HAS_WRITTEN_DP: OUT STD_LOGIC;
	     --OUTPUT
	     UNDERFLOW: OUT STD_LOGIC;
	     MEM_A_ADDRESS, MEM_B_ADDRESS: OUT UNSIGNED(9 DOWNTO 0);
	     Y_SAT: OUT SIGNED(7 DOWNTO 0));
END DP;

ARCHITECTURE BEH OF DP IS

SIGNAL ADDRESS_SIG_MEM_A_WR, ADDRESS_SIG_MEM_B_WR, ADDRESS_SIG_MEM_A_RD: UNSIGNED(9 DOWNTO 0) := (OTHERS => '0');
SIGNAL Y: SIGNED (10 DOWNTO 0);
SIGNAL MEM_A_HAS_WRITTEN_SIG: STD_LOGIC := '0';

COMPONENT MEM_A_WR_COUNTER IS
	PORT(CLK, RST, EN, START: IN STD_LOGIC;
	ADDR: OUT UNSIGNED(9 DOWNTO 0);
	MEM_A_HAS_WRITTEN_M: OUT STD_LOGIC);
END COMPONENT;
	
COMPONENT MEM_B_WR_COUNTER IS
	PORT(CLK, RST, EN, DONE: IN STD_LOGIC;      
        ADDR: OUT UNSIGNED(9 DOWNTO 0));				 
END COMPONENT;

COMPONENT MEM_A_READ_COUNTER IS
	PORT(CLK, RST, EN: IN STD_LOGIC;
	ADDR_B: IN UNSIGNED(9 DOWNTO 0);   
	ADDR: OUT UNSIGNED(9 DOWNTO 0));
END COMPONENT;
	

COMPONENT FILTERING_FUNCTION IS
PORT(X : IN SIGNED (7 DOWNTO 0);
     inv: IN SIGNED;
     LD, SH: IN STD_LOGIC_VECTOR(2 downto 0);
     loc: IN NATURAL;
     CLOCK, RESET, D, RST_SUM : IN STD_LOGIC;
     Y : OUT SIGNED (10 DOWNTO 0));
END COMPONENT;

COMPONENT SATURATOR IS
	PORT(EN: IN STD_LOGIC;
	     inp: IN SIGNED (10 DOWNTO 0);
	     outp : OUT SIGNED (7 DOWNTO 0));     
END COMPONENT;


BEGIN

C0: MEM_A_WR_COUNTER PORT MAP(CLOCK, RESET, WR_A, START, ADDRESS_SIG_MEM_A_WR, MEM_A_HAS_WRITTEN_SIG); 

MEM_A_HAS_WRITTEN_DP  <=  MEM_A_HAS_WRITTEN_SIG WHEN (WR_A = '1') ELSE '0';

MEM_A_ADDRESS <= ADDRESS_SIG_MEM_A_WR WHEN WR_A = '1' ELSE
	     	 ADDRESS_SIG_MEM_A_RD;

UNDERFLOW <= '1' WHEN( ADDRESS_SIG_MEM_A_RD > ADDRESS_SIG_MEM_B_WR) ELSE
	     '0';

C1: MEM_A_READ_COUNTER PORT MAP(CLOCK, RESET, UPDATE_ADD, ADDRESS_SIG_MEM_B_WR , ADDRESS_SIG_MEM_A_RD);

C2: MEM_B_WR_COUNTER PORT MAP(CLOCK, RESET, WR_B, DONE, ADDRESS_SIG_MEM_B_WR);

FILTERING: FILTERING_FUNCTION PORT MAP(X, INV, LD, SH, N_SHIFT, CLOCK, RESET, D, RESET_SUM, Y);

SAT: SATURATOR PORT MAP(EN_SAT, Y, Y_SAT);

MEM_B_ADDRESS <= ADDRESS_SIG_MEM_B_WR;

END BEH;

	     
	     